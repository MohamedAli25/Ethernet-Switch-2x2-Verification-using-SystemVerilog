module Switch(
    input clk,
    input rstN,
    input [31:0] inDataA,
    input insopA,
    input ineopA,
    input [31:0] inDataB,
    input insopB,
    input ineopB,
    output [31:0] outputA,
    output outsopA,
    output outeopA,
    output [31:0] outDataB,
    output outsopB,
    output outeopB,
    output portAStall,
    output portBStall
);

endmodule